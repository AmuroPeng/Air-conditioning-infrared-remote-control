`timescale 1ns / 1ps
module hongwai(clk,rst,key_1,IR_out,IR_outt,led_out);
input clk;
input rst;
input key_1; //����
wire [34:0] IR_in_data35;
wire [32:0] IR_in_data32;
output IR_out;
output led_out; //��ȫ���һ��ָ�����led��һ��
output IR_outt;
// output IR_outt_rev;

reg led;
reg [34:0] data35;
reg [32:0] data32;
reg [32:0] data32temp;

parameter t_38k    = 12'd3289;//125MHz/38kHz
parameter t_38k_half = 12'd1644;
parameter t_9ms    = 21'd1125000;//125MHz*9ms
parameter t_4_5ms  = 20'd562500;
parameter t_13_5ms = 21'd1687500;
parameter t_20000us = 22'd2500000;
parameter t_20750us = 22'd2593750;
parameter t_750us = 17'd93750;
parameter t_450us = 16'd56250;
parameter t_1500us = 18'd187500;
parameter t_1200us = 18'd150000;
parameter t_2250us = 19'd281250;

// �������ϵĹ���YB0F2ң�����ı���Э��
// parameter t_38k    = 12'd3289;//125MHz/38kHz
// parameter t_38k_half = 12'd1644;
// parameter t_9ms    = 21'd1125000;//125MHz*9ms
// parameter t_4_5ms  = 20'd562500;
// parameter t_13_5ms = 21'd1687500;
// parameter t_20000us = 22'd2500000;
// parameter t_20750us = 22'd2575000;
// parameter t_750us = 17'd75000;
// parameter t_450us = 16'd75000;
// parameter t_1500us = 18'd200000;
// parameter t_1200us = 18'd150000;
// parameter t_2250us = 19'd275000;

//38k��Ƶ----------------------------------------------//
reg  [12:0] cnt1;
wire  clk_38k;
always @(posedge clk or negedge rst)
    begin
        if(rst)
            begin
                cnt1 <= 0;
            end
        else if(cnt1 == t_38k)
                begin
                    cnt1 <= 0;
                end
            else cnt1 <= cnt1 + 1;
    end
assign  clk_38k = (cnt1<t_38k_half)?0:1;
//38k��Ƶ----------------------------------------------//

//״̬������----------------------------------------------//

parameter  IDEL       = 3'D0;        //��ʼ��״̬���ȴ���������
parameter  START      = 3'D1;        //��ʼ������ʼ�� 
parameter  SEND_35    = 3'D2;        //����35λ������
parameter  CONNECT    = 3'D3;        //����������
parameter  SEND_32    = 3'D4;        //����32λ������
reg   [2:0]     state;
reg             start_en;//��ʼ_ʹ��
wire            start_over;//��ʼ���Ƿ��ͽ���
reg             zero_en;
wire            zero_over;//��Щ�ж��Ƿ�����ı�����Ȼ������always��������ֵ��û���޸�ֻ�������жϣ�����wire��û��ë��
reg             one_en;
wire            one_over;
reg             connect_en;
wire            connect_over;
reg             data35_over;
reg             data32_over;
reg             idel_flag;
// reg             kaiguan;

reg   [5:0]     i;//��¼����Ŀǰ��λ��

always @(posedge clk or negedge rst)
    begin
        if(rst)
            begin
                state <= IDEL;
                start_en <= 0;
                zero_en <= 0;
                one_en <= 0;
                connect_en <= 0;
                // sendover <= 0;
                // shiftdata <= 0; 
                i <= 6'd34; //��data35����
                // DATA <= 8'D0;
                // kaiguan <= 1;
            end                   
        else 
            begin
                case(state)
                    IDEL:
                        begin
                            start_en <= 0;
                            zero_en <= 0;
                            one_en <= 0;
                            connect_en <= 0;
                            data35_over <= 0;
                            data32_over <= 0;
                            i <= 6'd34;//��data35����
                            led <= 0;//Ϩ��һյС��
                            idel_flag <= 1;
                            if(key_1)//�ػ�
                                begin
                                    state <= START;    
                                    data35 <= 35'b10000010000100000000010000001010010;
                                    data32 <= 33'b000010000000010000000000000001100;
                                    idel_flag <= 0;
                                end
                            else 
                                begin
                                    if(data32temp != data32)//����һ��˵��û����ָ��룬��һ����˵����Ҫ���е��Ʋ������
                                        begin//����Ŷ���Ǽ�begin&end�ˣ�����֮���else�ϱ���debug����T_T
                                            data35 <= IR_in_data35;
                                            data32 <= IR_in_data32;
                                            state <= START;
                                            idel_flag <= 1;
                                        end
                                    else state <= IDEL;//ƽʱһֱ��IDEL״̬�����
                                end
                        end
                    START:  //������ʼ��
                        begin
                            if(start_over)    
                                begin                                         
                                    start_en <= 0;
                                    state <= SEND_35;    
                                end
                            else 
                                begin
                                    start_en <= 1;
                                    state <= START;     
                                end     
                        end
                    SEND_35:    //����35λ������
                        begin
                            if(data35_over)
                                begin  
                                    i <= 6'd32;    //��data32����
                                    one_en <= 0;
                                    zero_en <= 0;
                                    state <= CONNECT;
                                end
                            else 
                                begin
                                    if(zero_over||one_over)   //1bit���ͽ���
                                        begin
                                            if (i==0) //�Ƿ������һλ
                                                data35_over <= 1;
                                            i <= i - 1; //����һλ
                                            one_en <= 0;
                                            zero_en <= 0;
                                        end
                                    else if(data35[i]) one_en <= 1; 
                                    else if(!data35[i]) zero_en <= 1;
                                    // else 
                                    //     begin
                                    //         i <= i ;
                                    //         one_en <= one_en;
                                    //         zero_en <= zero_en;
                                    //     end  
                                end
                        end
                    CONNECT:  //����������
                        begin
                            if(connect_over)    
                                begin                                         
                                    connect_en <= 0;
                                    state <= SEND_32;   
                                end
                            else 
                                begin
                                    connect_en <= 1;
                                    state <= CONNECT;     
                                end     
                        end
                    SEND_32:    //����32λ������
                        begin
                            if(data32_over)
                                begin  
                                    i <= 6'd34;    //��data35����
                                    one_en <= 0;
                                    zero_en <= 0;
                                    data32temp <= data32;//�����ͺ��ֵ��¼��������IDEL״̬���Ͻ����ж�
                                    state <= IDEL;
                                end
                            else 
                                begin
                                    if(zero_over||one_over)   //1bit���ͽ���
                                        begin
                                            if (i==0) //�Ƿ������һλ
                                                data32_over <= 1;
                                            i <= i - 1; //����һλ
                                            one_en <= 0;
                                            zero_en <= 0;
                                            led <= 1;//����һյС��
                                        end
                                    else if(data32[i]) one_en <= 1; 
                                    else if(!data32[i]) zero_en <= 1;
                                    // else 
                                    //     begin
                                    //         i <= i ;
                                    //         one_en <= one_en;
                                    //         zero_en <= zero_en;
                                    //     end  
                                end
                        end
                    default: state <= IDEL;
                endcase
            end //end all cases
    end
//״̬������----------------------------------------------//


//----------------------------------------------//
//�����룬9ms�ز���4.5ms����
reg    [20:0]cnt2;//@@@���ݳ��Ⱥ�13.5msһ��
wire         start_flag;
always @(posedge clk or negedge rst)
    begin
        if(rst)
            begin
                cnt2 <= 0;
            end
        else if(start_en)
                begin
                    if(cnt2 >= t_13_5ms)  cnt2 <= t_13_5ms+1;        
                    else cnt2 <= cnt2 + 1;
                end
            else cnt2  <= 0;         
    end
assign start_over = (cnt2 == t_13_5ms)?1:0;    
assign start_flag = (start_en&&(cnt2 >= t_9ms))?1:0;

//�����룬 750us�ز� 20000us����
reg    [21:0]     cnt5;//@@@���ݳ��Ⱥ�20000usһ��
wire              finish_flag;
always @(posedge clk or negedge rst)
    begin
        if(rst)
            begin
                cnt5 <= 0;
            end
        else if(connect_en)
                begin
                    if(cnt5 >= t_20750us)  cnt5 <= t_20750us+1;        
                    else cnt5 <= cnt5 + 1;
                end
            else cnt5  <= 0;         
    end
assign connect_over = (cnt5 == t_20750us)?1:0;    
assign connect_flag = (connect_en&&(cnt5 >= t_750us))?1:0;

//----------------------------------------------//
//����0, 560us�ز� + 560us����
reg    [17:0]     cnt3;// @@@���ݳ��Ⱥ�1200usһ��
wire              zero_flag;
always @(posedge clk or negedge rst)
    begin
        if(rst)
            begin
                cnt3 <= 0;
            end
        else if(zero_en)
            begin
                if(cnt3 >= t_1200us)  cnt3 <= t_1200us+1;        
                else cnt3 <= cnt3 + 1;
            end
        else cnt3  <= 0;         
    end
assign zero_over = (cnt3 == t_1200us)?1:0;    
assign zero_flag = (zero_en&&(cnt3 >= t_750us))?1:0;
    
//----------------------------------------------//
//����1, 560us�ز� + 1.68ms����
reg    [18:0]     cnt4;// @@@���ݳ��Ⱥ�t_2250usһ��
wire              one_flag;
always @(posedge clk or negedge rst)
    begin
        if(rst)
            begin
                cnt4 <= 0;
            end
        else if(one_en)
            begin
                if(cnt4 >= t_2250us)  cnt4 <= t_2250us+1;        
                else cnt4 <= cnt4 + 1;
            end
        else cnt4  <= 0;         
    end
assign one_over = (cnt4 == t_2250us)?1:0;    
assign one_flag = (one_en&&(cnt4 >= t_750us))?1:0;
    
wire   ir_out;
wire  IR_outt_rev;
assign ir_out = start_flag||zero_flag||one_flag||connect_flag||idel_flag;
assign IR_out = ir_out;
// assign IR_outt_rev = ~IR_outt;
assign IR_outt = (~ir_out)&&clk_38k;//38k�ز����ڵ͵�ƽʱ�ŵ��ƣ�����Ҫ����ir_out�ķ�

assign led_out = led;

endmodule